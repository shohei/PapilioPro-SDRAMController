module SDRAM_Controller (
	input clk,
	input reset,
	input [31:0] IO_Address,
	input [3:0] IO_Byte_Enable,
	input [31:0] IO_Write_Data,
	input IO_Addr_Strobe,
	input IO_Read_Strobe,
        output wire SDRAM_CLK,
        output wire SDRAM_CKE,
        output wire SDRAM_CS,
        output wire SDRAM_RAS,
        output wire SDRAM_CAS,
        output wire SDRAM_WE,
        output wire [1:0] SDRAM_DQM,
        output wire [12:0] SDRAM_ADDR,
        output wire [1:0] SDRAM_BA,
        inout [15:0] SDRAM_DATA,

	//output reg data_out_ready,
	//output reg cmd_ready,//MEMIORDY

        /* バス・インターフェース */
        input               WRMEM,  WRREG,
        output      [31:0]  RDATA0, RDATA1,
        output reg MEMIORDY,
        /* グラフィック表示回路 */
        input       [20:0]  DMEMADDR,
        /* キャプチャ回路 */
        //input       [23:1]  CMEMADDR,//22bit
        input       [20:0]  CMEMADDR,//22bit
        input       [15:0]  CMEMDOUT,
        input               CMEMnWE_asrt, CMEMnWE_deas,
        /* MODE信号のLED表示用 */
        output  reg [1:0]   MODE
);

   parameter sdram_address_width   = 22;
   parameter sdram_column_bits     =  8;
   parameter sdram_startup_cycles  = 14'd10100;//10100
   //parameter cycles_per_refresh  =  (64100*100)/4196-1;
   //parameter cycles_per_refresh  =  ((64100*100)/4196-1)/10;
   parameter cycles_per_refresh  =  770;//for 50MHz
   parameter start_of_col = 1'b0;
   parameter end_of_col = sdram_column_bits-2; //6
   parameter start_of_bank = sdram_column_bits-1; //7
   parameter end_of_bank   = sdram_column_bits; //6
   parameter start_of_row  = sdram_column_bits+1; //9
   parameter end_of_row    = sdram_address_width-2; //20
   parameter prefresh_cmd  = 10;

   wire [sdram_address_width-2:0] cmd_address;//20:0 //21bit
   assign cmd_address = IO_Address[sdram_address_width-2:0];//22-2:0=20:0 lower 21bit
   wire [3:0] cmd_byte_enable;
   assign cmd_byte_enable = IO_Byte_Enable;
   //assign cmd_byte_enable = 4'b0011;
   wire [31:0] cmd_data_in;
   assign cmd_data_in = IO_Write_Data;
   reg [31:0] data_out;
   assign RDATA0 = data_out;
   reg data_out_ready;//not using

   //assign MEMIORDY = (state==s_idle_in_1) ? 1'b1: 1'b0;
   always @(posedge clk) begin
        if(reset)
        	MEMIORDY <= 1'b0;
        else if(state==s_idle_in_1)
        	MEMIORDY <= 1'b1;
        else if(state==s_idle)
        	MEMIORDY <= 1'b0;//on for 2 clock(coz it's double clk speed)
   end
   
   //From page 37 of MT48LC16M16A2 datasheet
   //Name (Function)       CS# RAS# CAS# WE# DQM  Addr    Data
   //COMMAND INHIBIT (NOP)  H   X    X    X   X     X       X
   //NO OPERATION (NOP)     L   H    H    H   X     X       X
   //ACTIVE                 L   L    H    H   X  Bank/row   X
   //READ                   L   H    L    H  L/H Bank/col   X
   //WRITE                  L   H    L    L  L/H Bank/col Valid
   //BURST TERMINATE        L   H    H    L   X     X     Active
   //PRECHARGE              L   L    H    L   X   Code      X
   //AUTO REFRESH           L   L    L    H   X     X       X 
   //LOAD MODE REGISTER     L   L    L    L   X  Op-code    X 
   //Write enable           X   X    X    X   L     X     Active
   //Write inhibit          X   X    X    X   H     X     High-Z

   // Here are the commands mapped to constants   
   parameter CMD_UNSELECTED     =  4'b1000;
   parameter  CMD_NOP 		=  4'b0111;
   parameter  CMD_ACTIVE        =  4'b0011;
   parameter  CMD_READ          =  4'b0101;
   parameter  CMD_WRITE         =  4'b0100;
   parameter  CMD_TERMINATE     =  4'b0110;
   parameter  CMD_PRECHARGE     =  4'b0010;
   parameter  CMD_REFRESH       =  4'b0001;
   parameter  CMD_LOAD_MODE_REG =  4'b0000;

   parameter MODE_REG = 13'b0_0000_0010_0001;

   //wire cmd_enable = 1'b1;
   reg cmd_enable;
   always @(posedge clk) begin
      if(reset)
   	   cmd_enable <= 1'b0;
      else if(IO_Addr_Strobe)
   	   cmd_enable <= 1'b1;
      else if(state==s_open_in_1)
   	   cmd_enable <= 1'b0;
   end

   reg cmd_wr;

   reg [3:0] iob_command = CMD_NOP;
   reg [12:0] iob_address = 13'b0;
   reg [15:0] iob_data = 16'b0;
   reg [1:0] iob_dqm; 
   reg iob_cke = 1'b0;
   reg [1:0] iob_bank = 2'b0; 
   
   reg [15:0] iob_data_next      = 16'b0;
   reg [15:0] captured_data      = 16'b0;
   reg [15:0] captured_data_last = 16'b0;
   wire [15:0] sdram_din;
   
   parameter s_startup    = 5'd1,    
             s_idle_in_6  = 5'd2,
	     s_idle_in_5  = 5'd3,
	     s_idle_in_4  = 5'd4,
	     s_idle_in_3  = 5'd5,
	     s_idle_in_2  = 5'd6,
	     s_idle_in_1  = 5'd7,
             s_idle       = 5'd8,
             s_open_in_2  = 5'd9,
	     s_open_in_1  = 5'd10,
             s_write_1    = 5'd11,   
	     s_write_2    = 5'd12, 
	     s_write_3    = 5'd13, 
             s_read_1     = 5'd14, 
	     s_read_2     = 5'd15,
	     s_read_3     = 5'd16,
	     s_read_4     = 5'd17,
             s_precharge  = 5'd18;

   reg [4:0] state = s_startup;
   
   parameter [13:0] startup_refresh_max =14'b11_1111_1111_1111;//14'd16383
   reg [13:0] startup_refresh_count;

   // Indicate the need to refresh when the counter is 2048,
   // Force a refresh when the counter is 4096 - (if a refresh is forced, 
   // multiple refresshes will be forced until the counter is below 2048
   wire pending_refresh; 
   wire forcing_refresh; 
   assign pending_refresh = startup_refresh_count[11];
   assign forcing_refresh = startup_refresh_count[12];

   wire [12:0] addr_row;
   wire [12:0] addr_col;
   wire [1:0] addr_bank; 

   reg [3:0] dqm_sr = 4'b1111;
   
   reg save_wr = 1'b0;        
   reg [12:0] save_row;
   reg [1:0] save_bank;
   reg [12:0] save_col;
   reg [31:0] save_data_in;
   reg [3:0] save_byte_enable;
   
   reg ready_for_new = 1'b0;  
   reg got_transaction = 1'b0;
   
   reg can_back_to_back = 1'b0;

   reg iob_dq_hiz = 1'b1;

   reg [3:0] data_ready_delay;
   
  

   //tell the outside world when we can accept a new transaction;
   assign cmd_ready = ready_for_new;
   //----------------------------------------------------------------------------
   //-- Seperate the address into row / bank / address
   //----------------------------------------------------------------------------
   //parameter end_of_col = sdram_column_bits-2; //6
   //parameter start_of_bank = sdram_column_bits-1; //7
   //parameter end_of_bank   = sdram_column_bits; //6
   //parameter start_of_row  = sdram_column_bits+1; //9
   //parameter end_of_row    = sdram_address_width-2; //20
   //parameter prefresh_cmd  = 10;
   //parameter start_of_col = 1'b0;
   //parameter end_of_col = sdram_column_bits-2; //6
   //assign addr_row[end_of_row-start_of_row:0] = cmd_address[end_of_row:start_of_row];  //-- 12:0 <=  22:10 //11:0, 20:9, 12bit
   assign addr_row = {1'b0,cmd_address[end_of_row:start_of_row]};  //-- 12:0 <=  22:10 //11:0, 20:9, 12bit
   //assign addr_col[sdram_column_bits-1:0] = {cmd_address[end_of_col:start_of_col],1'b0}; // -- 8:0  <=  7:0 & '0' //7:0 ->{6:0},0
   assign addr_col = {5'b00000,cmd_address[end_of_col:start_of_col],1'b0}; // -- 8:0  <=  7:0 & '0' //7:0 ->{6:0},0
   assign addr_bank = cmd_address[end_of_bank:start_of_bank];//      -- 1:0  <=  9:8

   //-----------------------------------------------------------
   //-- Forward the SDRAM clock to the SDRAM chip - 180 degress 
   //-- out of phase with the control signals (ensuring setup and holdup 
  //----------------------------------------------------------
ODDR2 #(
	   .DDR_ALIGNMENT("NONE"),
	   .INIT(1'b0), 
	   .SRTYPE("SYNC")
   )
   ODDR_inst (
	   .Q(SDRAM_CLK),
	   .C0(clk),
           .C1(~clk),
	   .CE(1'b1), 
	   .R(1'b0), 
	   .S(1'b0), 
	   .D0(1'b0), 
	   .D1(1'b1)
   );

   //j-----------------------------------------------
   //j--!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
   //j--!! Ensure that all outputs are registered. !!
   //j--!! Check the pinout report to be sure      !!
   //j--!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
   //j-----------------------------------------------
   assign SDRAM_CKE = iob_cke;
   assign SDRAM_CS = iob_command[3];
   assign SDRAM_RAS = iob_command[2];
   assign SDRAM_CAS = iob_command[1];
   assign SDRAM_WE = iob_command[0];
   assign SDRAM_DQM = iob_dqm;
   assign SDRAM_BA = iob_bank;
   assign SDRAM_ADDR = iob_address;
   
   //---------------------------------------------------------------
   //-- Explicitly set up the tristate I/O buffers on the DQ signals
   //---------------------------------------------------------------
genvar i;
generate
for(i=0;i<16;i=i+1)
    begin
    IOBUF #(
    	.DRIVE(12),
    	.IOSTANDARD("LVTTL"),
    	.SLEW("FAST")
           )
         IOBUF_inst(
    	     .O (sdram_din[i]),
    	     .IO(SDRAM_DATA[i]), 
    	     .I (iob_data[i]), 
    	     .T (iob_dq_hiz)
         );
    end
endgenerate


always @(posedge clk) begin
   if(reset)
	   cmd_wr <= 1'b0;
   else if(WRMEM)
	   cmd_wr <= 1'b1;
   else if(state==s_write_2)
	   cmd_wr <= 1'b0;
end
                                     
always @(posedge clk) begin
         captured_data  <= sdram_din;
end

always @(posedge clk) begin
         captured_data_last <= captured_data;
         //------------------------------------------------
         //-- countdown for initialisation & refresh
         //------------------------------------------------
	 if(reset)
		startup_refresh_count <= startup_refresh_max-sdram_startup_cycles;//16383-10100=6283
	 else
                startup_refresh_count <= startup_refresh_count+14'd1;
         //-------------------------------------------------------------------
         //-- It we are ready for a new tranasction and one is being presented
         //-- then accept it. Also remember what we are reading or writing,
         //-- and if it can be back-to-backed with the last transaction
         //-------------------------------------------------------------------
	 if (ready_for_new==1'b1 && cmd_enable==1'b1) begin
	    if(save_bank==addr_bank&&save_row==addr_row)
               can_back_to_back <= 1'b1;
            else 
               can_back_to_back <= 1'b0;
            
            save_row         <= addr_row;
            save_bank        <= addr_bank;
            save_col         <= addr_col;
            save_wr          <= cmd_wr; 
            save_data_in     <= cmd_data_in;
            save_byte_enable <= cmd_byte_enable;
            got_transaction  <= 1'b1;
            ready_for_new    <= 1'b0;
         end
         //------------------------------------------------
         //-- Handle the data coming back from the 
         //-- SDRAM for the Read transaction
         //------------------------------------------------
         data_out_ready <= 1'b0;
	 if (data_ready_delay[0]==1'b1) begin
            data_out       <= {captured_data,captured_data_last};
            //data_out       <= {captured_data_last,captured_data};
            data_out_ready <= 1'b1;
         end
         //----------------------------------------------------------------------------
         //-- update shift registers used to choose when to present data to/from memory
         //----------------------------------------------------------------------------
         data_ready_delay <= {1'b0,data_ready_delay[3:1]};
         iob_dqm          <= dqm_sr[1:0]; //lower 2bit
         dqm_sr           <= {2'b11,dqm_sr[3:2]};//upper 2bit

         case (state)
	     s_startup: begin
               //------------------------------------------------------------------------
               //-- This is the initial startup state, where we wait for at least 100us
               //-- before starting the start sequence
               //-- 
               //-- The initialisation is sequence is 
               //--  * de-assert SDRAM_CKE
               //--  * 100us wait, 
               //--  * assert SDRAM_CKE
               //--  * wait at least one cycle, 
               //--  * PRECHARGE
               //--  * wait 2 cycles
               //--  * REFRESH, 
               //--  * tREF wait
               //--  * REFRESH, 
               //--  * tREF wait 
               //--  * LOAD_MODE_REG 
               //--  * 2 cycles wait
               //------------------------------------------------------------------------
               iob_cke <= 1'b1;
               
               //-- All the commands during the startup are NOPS, except these
	       
               //max = 16383
	       if (startup_refresh_count == startup_refresh_max-14'd31) begin //16352
                  //-- ensure all rows are closed
                  iob_command     <= CMD_PRECHARGE;
                  iob_address[prefresh_cmd] <= 1'b1; // -- all banks
                  iob_bank    <= 2'b0;
	       end
               else if (startup_refresh_count == startup_refresh_max-14'd23)//16360
                  //-- these refreshes need to be at least tREF (66ns) apart
                  iob_command     <= CMD_REFRESH;
               else if (startup_refresh_count == startup_refresh_max-14'd15)//16368
                  iob_command     <= CMD_REFRESH;
	       else if (startup_refresh_count == startup_refresh_max-14'd7) begin //16376-- Now load the mode register
                       iob_command     <= CMD_LOAD_MODE_REG;
                       iob_address     <= MODE_REG;
	       end
               //------------------------------------------------------
               //-- if startup is coomplete then go into idle mode,
               //-- get prepared to accept a new command, and schedule
               //-- the first refresh cycle
               //------------------------------------------------------
	       if (startup_refresh_count == 14'd0) begin
                  state           <= s_idle;
                  ready_for_new   <= 1'b1;
                  got_transaction <= 1'b0;
                  startup_refresh_count <= 14'd2048 - cycles_per_refresh+14'd1;
		  iob_command <= CMD_NOP;
	       end
               
               
            end
            s_idle_in_6 : state <= s_idle_in_5;
            s_idle_in_5 : state <= s_idle_in_4;
            s_idle_in_4 : state <= s_idle_in_3;
            s_idle_in_3 : state <= s_idle_in_2;
            s_idle_in_2 : state <= s_idle_in_1;
	    s_idle_in_1 : begin
		    state <= s_idle;
		    iob_command <= CMD_NOP;
	    end

	    s_idle : begin
               //-- Priority is to issue a refresh if one is outstanding
	       if (pending_refresh == 1'b1 || forcing_refresh == 1'b1) begin
                  //------------------------------------------------------------------------
                  //-- Start the refresh cycle. 
                  //-- This tasks tRFC (66ns), so 6 idle cycles are needed @ 100MHz
                  //------------------------------------------------------------------------
                  state       <= s_idle_in_6;
                  iob_command <= CMD_REFRESH;
                  startup_refresh_count <= startup_refresh_count - cycles_per_refresh+1;//
	       end
	       else if (got_transaction == 1'b1) begin
                  //--------------------------------
                  //-- Start the read or write cycle. 
                  //-- First task is to open the row
                  //--------------------------------
                  state       <= s_open_in_2;
                  iob_command <= CMD_ACTIVE;
                  iob_address <= save_row;
                  iob_bank    <= save_bank;
               end 

	    end
            //--------------------------------------------
            //-- Opening the row ready for reads or writes
            //--------------------------------------------
	    s_open_in_2 : begin
	      state <= s_open_in_1;
              //iob_dq_hiz  <= 1'b0;//open IO buffer: though this not be all-right for reading...
      	    end

	    s_open_in_1 : begin
               //-- still waiting for row to open
	       if (save_wr == 1'b1) begin
                  state       <= s_write_1;
                  iob_dq_hiz  <= 1'b0;
                  iob_data    <= save_data_in[15:0];// -- get the DQ bus out of HiZ early
	       end
	       else begin
                  iob_dq_hiz  <= 1'b1;
                  state       <= s_read_1;
	       end
               //-- we will be ready for a new transaction next cycle!
               ready_for_new   <= 1'b1; 
               got_transaction <= 1'b0;                  
              end

            //----------------------------------
            //-- Processing the read transaction
            //----------------------------------
	    s_read_1 : begin
               state           <= s_read_2;
               iob_command     <= CMD_READ;
               iob_address     <= save_col; 
               iob_bank        <= save_bank;
               iob_address[prefresh_cmd] <= 1'b0; //-- A10 actually matters - it selects auto precharge
               
               //-- Schedule reading the data values off the bus
               data_ready_delay[3]   <= 1'b1;
               
               //-- Set the data masks to read all bytes
               iob_dqm  <= 2'b0;
               dqm_sr[1:0] <= 2'b0;
               
            end
	    s_read_2 : begin
               state <= s_read_3;
               if (forcing_refresh == 1'b0 && got_transaction == 1'b1 && can_back_to_back == 1'b1) begin
		 if (save_wr == 1'b0) begin
                     state           <= s_read_1;
                     ready_for_new   <= 1'b1;// -- we will be ready for a new transaction next cycle!
                     got_transaction <= 1'b0;
	         end
	       end 
            end
	    s_read_3 : begin
               state <= s_read_4;
               if (forcing_refresh == 1'b0 && got_transaction == 1'b1 && can_back_to_back == 1'b1) begin
		   if (save_wr == 1'b0) begin
                     state           <= s_read_1;
                     ready_for_new   <= 1'b1;// -- we will be ready for a new transaction next cycle!
                     got_transaction <= 1'b0;
	           end
	       end

            end
	    s_read_4 : begin
               state <= s_precharge;
               //-- can we do back-to-back read?
	       if (forcing_refresh == 1'b0 && got_transaction == 1'b1 && can_back_to_back == 1'b1)  begin
		 if (save_wr == 1'b0) begin
                     state           <= s_read_1;
                     ready_for_new   <= 1'b1; //-- we will be ready for a new transaction next cycle!
                     got_transaction <= 1'b0;
	          end
                  else
                     state <= s_open_in_2; //-- we have to wait for the read data to come back before we swutch the bus into HiZ
               end
	    end
            //------------------------------------------------------------------
            //-- Processing the write transaction
            //-------------------------------------------------------------------
	    s_write_1 : begin
               state              <= s_write_2;
               iob_command        <= CMD_WRITE;
               iob_address        <= save_col; 
               iob_address[prefresh_cmd]    <= 1'b0; //-- A10 actually matters - it selects auto precharge
               iob_bank           <= save_bank;
               iob_dqm            <= ~save_byte_enable[1:0];    
               dqm_sr[1:0] <= ~save_byte_enable[3:2];    
               iob_data           <= save_data_in[15:0];
               iob_data_next      <= save_data_in[31:16];
               
            end
	    s_write_2 : begin
               state           <= s_write_3;
               iob_data        <= iob_data_next; //comment out for debug
               //dqm_sr[1:0] <= ~save_byte_enable[1:0]; //debug
               //-- can we do a back-to-back write?
	       if (forcing_refresh == 1'b0 && got_transaction == 1'b1 && can_back_to_back == 1'b1)begin
		 if (save_wr == 1'b1) begin
                     //-- back-to-back write?
                     state           <= s_write_1;
                     ready_for_new   <= 1'b1;
                     got_transaction <= 1'b0;
                  //-- Although it looks right in simulation you can't go write-to-read 
                  //-- here due to bus contention, as iob_dq_hiz takes a few ns.
		  end
	       end
         
            end
	    s_write_3 : begin// must wait tRDL, hence the extra idle state
               //-- back to back transaction?
	       if (forcing_refresh == 1'b0 && got_transaction == 1'b1 && can_back_to_back == 1'b1) begin
		  if (save_wr == 1'b1) begin
                     //-- back-to-back write?
                     state           <= s_write_1;
                     ready_for_new   <= 1'b1;
                     got_transaction <= 1'b0;
	          end
		  else begin
                     //-- write-to-read switch?
                     state           <= s_read_1;
                     iob_dq_hiz      <= 1'b1;
                     ready_for_new   <= 1'b1; //-- we will be ready for a new transaction next cycle!
                     got_transaction <= 1'b0;                  
	          end
	       end
	       else begin
                    iob_dq_hiz         <= 1'b1;//comment out for debug
		    //iob_data <= save_data_in[31:16];//debug
		    iob_data <= save_data_in[15:0];//debug
		    //iob_command <= CMD_TERMINATE;
                    state              <= s_precharge;
	       end //else
            end //s_write_3
            //-------------------------------------------------------------------
            //-- Closing the row off (this closes all banks)
            //-------------------------------------------------------------------
	    s_precharge : begin
	       iob_dq_hiz <= 1'b1;//debug
               state           <= s_idle_in_3;
               iob_command     <= CMD_PRECHARGE;
               iob_address[prefresh_cmd] <= 1'b1; //-- A10 actually matters - it selects all banks or just one
            end

            //-------------------------------------------------------------------
            //-- We should never get here, but if we do then reset the memory
            //-------------------------------------------------------------------
	    default : begin
               state                 <= s_startup;
               ready_for_new         <= 1'b0;
               startup_refresh_count <= startup_refresh_max-sdram_startup_cycles; //14bit
            end
         endcase

	 if (reset) begin //-- Sync reset 
            state                 <= s_startup;
            ready_for_new         <= 1'b0;
            startup_refresh_count <= startup_refresh_max-sdram_startup_cycles; //14bit
         end

end


/* メモリアクセス・モード設定レジスタ */
parameter DISPMODE=2'b00, CAPTMODE=2'b01, MCSMODE=2'b10;

always @( posedge clk) begin
    if ( reset )
        MODE <= 2'h0;
    else if ( WRREG & IO_Byte_Enable[0] )
        MODE <= IO_Write_Data[1:0];
end

/* メモリ読み出し信号 */
wire RDMEM = (IO_Address[31:24]==8'hc0) & IO_Read_Strobe;

/* MCSモード時のメモリ信号 */
//reg  [23:1]  MMEMADDR;
reg  [20:0]  MMEMADDR; //21bit address from MCS or other buses
reg          MMEMnOE, MMEMnWE, MMEMnUB, MMEMnLB;

reg         MEMnOE, MEMnWE, MEMnUB, MEMnLB;

/*TODO: メモリ信号切り替え */
/*
always @* begin
    case ( MODE )
        DISPMODE:   begin
			SDRAM_BA <= DMEMADDR[20:19];
                        SDRAM_ADDR[11:0] <= DMEMADDR[19:7]; //12 bit ROW ADDRESS(for lower 16bit data)
                        //SDRAM_ADDR[7:0] = {DMEMADDR[6:0],1'b0}; //8 bit COL ADDRESS(for lower 16bit data)
                        MEMnOE  = 1'b0; //VGA read from SDRAM
                        MEMnUB  = 1'b0;
                        MEMnLB  = 1'b0;
                    end
        CAPTMODE:   begin
			SDRAM_BA <= CMEMADDR[20:19];
                        SDRAM_ADDR <= CMEMADDR;
                        //SDRAM_ADDR[7:0] = {CMEMADDR[6:0],1'b0}; //8 bit COL ADDRESS(for lower 16bit data)
                        MEMnOE  = 1'b1; //CAMERA write to SDRAM
                        MEMnUB  = 1'b0;
                        MEMnLB  = 1'b0;
                    end
        MCSMODE:    begin
                        MEMnOE  = MMEMnOE; //read or write from MCS
                        MEMnUB  = MMEMnUB;
                        MEMnLB  = MMEMnLB;
                    end
        default:    begin
                        SDRAM_BA <= 2'b0;
                        SDRAM_ADDR <= 12'b0;
                        MEMnOE  = 1'b1;
                        MEMnUB  = 1'b1;
                        MEMnLB  = 1'b1;
                    end
    endcase
end
*/

endmodule

